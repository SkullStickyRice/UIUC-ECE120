-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION vending_machine_struct_config OF vending_machine IS
   FOR struct
   END FOR;
END vending_machine_struct_config;
